../../halfband_polyphase_test.srcs/sources_1/new/halfband_polyphase_fir.sv